// Blink an LED provided an input clock
/* module */
module top (hwclk, led1, led2, led3, led4, led5);
    /* I/O */
    input hwclk;
    output led1;
    output led2;
    output led3;
    output led4;
    output led5;

endmodule
